module fetch (
    
);

endmodule